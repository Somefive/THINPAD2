----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:07:08 11/17/2016 
-- Design Name: 
-- Module Name:    RamBlock - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity RamBlock is
    Port ( RegX : in STD_LOGIC_VECTOR (15 downto 0);
			  RegY : in STD_LOGIC_VECTOR (15 downto 0);
			  ALU : in STD_LOGIC_VECTOR(15 downto 0);
			  PC : in STD_LOGIC_VECTOR(15 downto 0);
			  RamControl : in STD_LOGIC_VECTOR(2 downto 0);
			  Finish : out STD_LOGIC;
			  Output : out STD_LOGIC_VECTOR(15 downto 0);
			  Ins : out STD_LOGIC_VECTOR(15 downto 0);
			  RAM1ADDR : out  STD_LOGIC_VECTOR (17 downto 0);
           RAM1DATA : inout  STD_LOGIC_VECTOR (15 downto 0);
           RAM1_EN : out  STD_LOGIC;
           RAM1_OE : out  STD_LOGIC;
           RAM1_WE : out  STD_LOGIC;
			  RAM2ADDR : out  STD_LOGIC_VECTOR (17 downto 0);
           RAM2DATA : inout  STD_LOGIC_VECTOR (15 downto 0);
           RAM2_EN : out  STD_LOGIC;
           RAM2_OE : out  STD_LOGIC;
           RAM2_WE : out  STD_LOGIC;
			  DATA_READY : in  STD_LOGIC;
           RDN : out  STD_LOGIC;
           TBRE : in  STD_LOGIC;
           TSRE : in  STD_LOGIC;
           WRN : out  STD_LOGIC;
           CLK : in  STD_LOGIC);
end RamBlock;

architecture Behavioral of RamBlock is
signal state: integer range 0 to 7:=0;
begin
	
	RAM1_EN <= '1';
	RAM1_OE <= '1';
	RAM1_WE <= '1';
	RAM2_EN <= '0';
	
	process(RamControl,CLK)
	begin
		if(CLK'event and CLK='1')then
			case RamControl is
				when "001" => -- Read Ins
					RAM2ADDR <= "00"&PC;
					RAM2DATA <= (others => 'Z');
					RAM2_OE <= '0';
					FINISH <= '0';
				when "011" => -- Finish Read Ins
					Ins <= RAM2DATA;
					RAM2_OE <= '1';
				when "010" => -- Read Data
					if(ALU(15 downto 1)="110111110000000")then
						RAM1DATA <= (others => 'Z');
						RDN <= '1';
						state <= 1;
					else
						RAM2ADDR <= "00"&ALU;
						RAM2DATA <= (others => 'Z');
						RAM2_OE <= '0';
						state <= 0;
					end if;
					FINISH <= '0';
				when "100" => -- Finish Read Data
					case state is
						when 0 =>
							Output <= RAM2DATA;
							RDN <= '1';
							FINISH <= '1';
						when 1 =>
							if(DATA_READY='0')then
								RDN<='1';
								RAM1DATA <= (others => 'Z');
							else
								RDN<='0';
								state <= 2;
							end if;
						when 2 =>
							Output <= "00000000"&RAM1DATA(7 downto 0);
							RDN<='1';
							FINISH<='1';
						when others =>
					end case;
				when "101" => --Write RegX
					if(ALU(15 downto 1)="110111110000000")then
						if(ALU(0)='0')then
							RAM1DATA <= RegX;
						else
							RAM1DATA <= "000000000000000"&DATA_READY;
						end if;
						WRN <= '0';
						state <= 1;
					else
						RAM2ADDR <= "00"&ALU;
						RAM2DATA <= RegX;
						RAM2_WE <= '0';
						state <= 0;
					end if;
				when "110" => --Write RegY
					if(ALU(15 downto 1)="110111110000000")then
						if(ALU(0)='0')then
							RAM1DATA <= RegY;
						else
							RAM1DATA <= "000000000000000"&DATA_READY;
						end if;
						WRN <= '0';
						state <= 1;
					else
						RAM2ADDR <= "00"&ALU;
						RAM2DATA <= RegY;
						RAM2_WE <= '0';
						state <= 0;
					end if;
				when "111" => --Finish Write Reg
					case state is
						when 0 =>
							WRN <= '1';
							RAM2_WE <= '1';
							FINISH <= '1';
						when 1 =>
							WRN <= '1';
							if(TBRE='1')then
								state <= 2;
							end if;
						when 2 =>
							if(TSRE='1')then
								state <= 0;
							end if;
						when others =>
					end case;
				when others =>
					RAM2_WE <= '1';
					RAM2_OE <= '1';
					WRN <= '1';
					RDN <= '1';
					FINISH <= '0';
			end case;
		end if;
	end process;

end Behavioral;

